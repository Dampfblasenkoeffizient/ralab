-- Clara Heilig