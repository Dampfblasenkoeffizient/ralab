library ieee;
use ieee.std_logic_1164.all;

--use work.constant_package.all;


entity my_alu is generic(
        G_DATA_WIDTH_GEN : integer := 32;
        G_ALU_OPCODE_WIDTH : integer := 4
    ); 
    port(
        pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
        pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
        pi_opcode    : in  std_logic_vector(G_ALU_OPCODE_WIDTH - 1 downto 0);
        po_result    : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
        po_carryOut  : out std_logic
    );
end my_alu;

architecture my_alu_arch of my_alu is
--    component and_alu
--            pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--            pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--            po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0)
--        );
--    end component;
--    component or_alu
--        port(
--            pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--            pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--            po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0)
--        );
--    end component;
--    component xor_alu
--        port(
--            pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--            pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--            po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0)
--        );
--    end component;
--    component sll_alu
--    port(
--        pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0)
--    );
--    end component;
--    component srl_alu
--    port(
--        pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0)
--    );
--    end component;
--    component sra_alu
--    port(
--        pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0)
--    );
--    end component;
--    component add_alu
--    port(
--        pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        po_carry     : out std_logic
--    );
--    end component;
--    component sub_alu
--    port(
--        pi_opa       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        pi_opb       : in  std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        po_out       : out std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
--        po_carry     : out std_logic
--    );
--    end component;

    signal s_and_result : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_or_result  : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_xor_result : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_sll_result : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_srl_result : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_sra_result : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_add_result : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_sub_result : std_logic_vector(G_DATA_WIDTH_GEN - 1 downto 0);
    signal s_carry : std_logic;
    
    begin

    and_alu_inst : entity work.and_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_and_result);
    or_alu_inst  : entity work.or_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_or_result);
    xor_alu_inst : entity work.xor_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_xor_result);
    sll_alu_inst : entity work.sll_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_sll_result);
    srl_alu_inst : entity work.srl_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_srl_result);
    sra_alu_inst : entity work.sra_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_sra_result);
    add_alu_inst : entity work.add_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_add_result, s_carry);
    sub_alu_inst : entity work.sub_alu generic map(G_DATA_WIDTH_GEN) port map(pi_opa, pi_opb, s_sub_result, s_carry);

        process(pi_opcode)
        variable v_opcode : std_logic_vector(G_ALU_OPCODE_WIDTH - 1 downto 0) := pi_opcode; --not static enough :( 
        begin 
            case v_opcode is
                when AND_ALU_OP => po_result <= s_and_result;
                when OR_ALU_OP => po_result <= s_or_result;
                when XOR_ALU_OP => po_result <= s_xor_result;
                when SLL_ALU_OP => po_result <= s_sll_result;
                when SRL_ALU_OP => po_result <= s_srl_result;
                when SRA_ALU_OP => po_result <= s_sra_result;
                when ADD_ALU_OP => po_result <= s_add_result;
                when SUB_ALU_OP => po_result <= s_sub_result;
                when others => po_result <= (others => '0');
            end case;
            po_carryOut <= s_carry;
        end process;
end architecture my_alu_arch;
    